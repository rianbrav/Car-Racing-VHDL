library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ram_catodo is
	port(data: in std_logic_vector(7 downto 0);
	add: in std_logic_vector(6 downto 0);
	modo: in std_logic;
	q: out std_logic_vector(7 downto 0));
end ram_catodo;
architecture sol of ram_catodo is
begin
		process(modo,add)
			begin
				if modo='1' then 
					case add is
					   when "0000000" => q<="00000000";
						when "0000001" => q<="00000000";----cuadro1
						when "0000010" => q<="10000000";
						when "0000011" => q<="00000010";----cuadro1
						when "0000100" => q<="00000000";----cuadro2
						when "0000101" => q<="10000000";
						when "0000110" => q<="00000010";
						when "0000111" => q<="00100000";----cuadro2
						when "0001000" => q<="00000000";----cuadro3
						when "0001001" => q<="10000000";
						when "0001010" => q<="00000010";
						when "0001011" => q<="00100000";
						when "0001100" => q<="00001000";---cuadro3
						when "0001101" => q<="00000000";---cuadro4
						when "0001110" => q<="10000000";
						when "0001111" => q<="00000010";
						when "0010000" => q<="00100000";
						when "0010001" => q<="00001000";---cuadro4
						when "0010010" => q<="10000000";---cuadro5
						when "0010011" => q<="00000010";
						when "0010100" => q<="00100000";
						when "0010101" => q<="00001000";
						when "0010110" => q<="00000010";---cuadro5
						when "0010111" => q<="00000000";---cuadro6
						when "0011000" => q<="00000010";
						when "0011001" => q<="00100000";
						when "0011010" => q<="00001000";
						when "0011011" => q<="00000010";
						when "0011100" => q<="01000000";---cuadro6
						when "0011101" => q<="00000010";---cuadro7
						when "0011110" => q<="00100000";
						when "0011111" => q<="00001000";
						when "0100000" => q<="00000010";
						when "0100001" => q<="01000000";---cuadro7
						when "0100010" => q<="00000000";---cuadro8
						when "0100011" => q<="00100000";
						when "0100100" => q<="00001000";
						when "0100101" => q<="00000010";
						when "0100110" => q<="01000000";
						when "0100111" => q<="00010000";---cuadro8
						when "0101000" => q<="00100000";---cuadro9
						when "0101001" => q<="00001000";
						when "0101010" => q<="00000010";
						when "0101011" => q<="01000000";
						when "0101100" => q<="00010000";
						when "0101101" => q<="00000100";---cuadro9
						when "0101110" => q<="00001000";---cuadro10
						when "0101111" => q<="00000010";
						when "0110000" => q<="01000000";
						when "0110001" => q<="00010000";
						when "0110010" => q<="00000100";---cuadro10
						when "0110011" => q<="00000000";---cuadro11
						when "0110100" => q<="00000010";
						when "0110101" => q<="01000000";
						when "0110110" => q<="00010000";
						when "0110111" => q<="00000100";
						when "0111000" => q<="00100000";---cuadro11
						when "0111001" => q<="00000010";---cuadro12
						when "0111010" => q<="01000000";
						when "0111011" => q<="00010000";
						when "0111100" => q<="00000100";
						when "0111101" => q<="00100000";
						when "0111110" => q<="00000001";---cuadro12
						when "0111111" => q<="01000000";---cuadro13
						when "1000000" => q<="00010000";
						when "1000001" => q<="00000100";
						when "1000010" => q<="00100000";
						when "1000011" => q<="00000001";
						when "1000100" => q<="01000000";---cuadro13
						when "1000101" => q<="00000000";---cuadro14
						when "1000110" => q<="00010000";
						when "1000111" => q<="00000100";
						when "1001000" => q<="00100000";
						when "1001001" => q<="00000001";
						when "1001010" => q<="01000000";
						when "1001011" => q<="00000100";---cuadro14
						when "1001100" => q<="00010000";---cuadro15
						when "1001101" => q<="00000100";
						when "1001110" => q<="00100000";
						when "1001111" => q<="00000001";
						when "1010000" => q<="01000000";
						when "1010001" => q<="00000100";---cuadro15
						when "1010010" => q<="00000100";---cuadro16
						when "1010011" => q<="00100000";
						when "1010100" => q<="00000001";
						when "1010101" => q<="01000000";
						when "1010110" => q<="00000100";
						when "1010111" => q<="10000000";---cuadro16
						when "1011000" => q<="00000000";---cuadro17
						when "1011001" => q<="00100000";
						when "1011010" => q<="00000001";
						when "1011011" => q<="01000000";
						when "1011100" => q<="00000100";
						when "1011101" => q<="10000000";
						when "1011110" => q<="00001000";---cuadro17
						when "1011111" => q<="00100000";---cuadro18
						when "1100000" => q<="00000001";
						when "1100001" => q<="01000000";
						when "1100010" => q<="00000100";
						when "1100011" => q<="10000000";
						when "1100100" => q<="00001000";
						when "1100101" => q<="01000000";---cuadro18
						when "1100110" => q<="00000001";---cuadro19
						when "1100111" => q<="01000000";
						when "1101000" => q<="00000100";
						when "1101001" => q<="10000000";
						when "1101010" => q<="00001000";
						when "1101011" => q<="01000000";
						when "1101100" => q<="00000010";---cuadro19
						when "1101101" => q<="01000000";---cuadro20
						when "1101110" => q<="00000100";
						when "1101111" => q<="10000000";
						when "1110000" => q<="00001000";
						when "1110001" => q<="01000000";
						when "1110010" => q<="00000010";---cuadro20
						when "1110011" => q<="00000100";---cuadro21
						when "1110100" => q<="10000000";
						when "1110101" => q<="00001000";
						when "1110110" => q<="01000000";
						when "1110111" => q<="00000010";
						when "1111000" => q<="00010000";---cuadro21
						when "1111001" => q<="00000000";---cuadro22
						when "1111010" => q<="10000000";
						when "1111011" => q<="00001000";
						when "1111100" => q<="01000000";
						when "1111101" => q<="00000010";
						when "1111110" => q<="00010000";
						when "1111111" => q<="01000000";
					end case;
				else
					q <= "00000000";
				end if;
	end process;
end sol;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ram_puntuaciones is
	port(data: in std_logic_vector(10 downto 0);
	add: in std_logic_vector(3 downto 0);
	modo_escritura: in std_logic;
   cambio_direccion: out std_logic;
   cambiar_estado: out std_logic;	
	q: out std_logic_vector(10 downto 0);
	salida: out std_logic_vector(10 downto 0));
end ram_puntuaciones;
architecture sol of ram_puntuaciones is
	signal r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15: std_logic_vector(10 downto 0):="00000000000";
	signal respaldo0, respaldo1, respaldo2, respaldo3, respaldo4, respaldo5, respaldo6, respaldo7, respaldo8, respaldo9, respaldo10, respaldo11, respaldo12, respaldo13, respaldo14, respaldo15: std_logic_vector(10 downto 0):="00000000000";
begin
	process(modo_escritura,add,data,respaldo0,respaldo1,respaldo2,respaldo3,respaldo4,respaldo5,respaldo6,respaldo7,respaldo8,respaldo9,respaldo10,respaldo11,respaldo12,respaldo13,respaldo14,r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15)
	begin
		q<="00000000000"; salida<="00000000000";
		if modo_escritura='1' then --escritura
			case add is
				when "0000" => if data > r0 then r0 <= data; end if;
									salida <= r0;
									cambio_direccion <= '1';
				when "0001" => if respaldo0 > r1 then r1 <= respaldo0;
									elsif data > r1 then r1 <= data; end if;
									salida <= r1;
									cambio_direccion <= '1';
				when "0010" => if respaldo0 > r2 then r2 <= respaldo0;
									elsif respaldo1 > r2 then r2 <= respaldo1;
									elsif data > r2 then r2 <= data; end if;
									salida <= r2;
									cambio_direccion <= '1'; 
				when "0011" => if respaldo0 > r3 then r3 <= respaldo0;
									elsif respaldo1 > r3 then r3 <= respaldo1;
									elsif respaldo2 > r3 then r3 <= respaldo2;
									elsif data > r3 then r3 <= data; end if;
									salida <= r3;
									cambio_direccion <= '1';
				when "0100" => if respaldo0 > r4 then r4 <= respaldo0;
									elsif respaldo1 > r4 then r4 <= respaldo1; 
									elsif respaldo2 > r4 then r4 <= respaldo2; 
									elsif respaldo3 > r4 then r4 <= respaldo3;
									elsif data > r4 then r4 <= data; end if;
									salida <= r4;
									cambio_direccion <= '1';
				when "0101" => if respaldo0 > r5 then r5 <= respaldo0;
									elsif respaldo1 > r5 then r5 <= respaldo1; 
									elsif respaldo2 > r5 then r5 <= respaldo2; 
									elsif respaldo3 > r5 then r5 <= respaldo3; 
									elsif respaldo4 > r5 then r5 <= respaldo4; 
									elsif data > r5 then r5 <= data; end if;
									salida <= r5;
									cambio_direccion <= '1';
				when "0110" => if respaldo0 > r6 then r6 <= respaldo0;
									elsif respaldo1 > r6 then r6 <= respaldo1;
									elsif respaldo2 > r6 then r6 <= respaldo2;
									elsif respaldo3 > r6 then r6 <= respaldo3;
									elsif respaldo4 > r6 then r6 <= respaldo4;
									elsif respaldo5 > r6 then r6 <= respaldo5;
									elsif data > r6 then r6 <= data; end if;
									salida <= r6;
									cambio_direccion <= '1';
				when "0111" => if respaldo0 > r7 then r7 <= respaldo0;
									elsif respaldo1 > r7 then r7 <= respaldo1;
									elsif respaldo2 > r7 then r7 <= respaldo2;
									elsif respaldo3 > r7 then r7 <= respaldo3;
									elsif respaldo4 > r7 then r7 <= respaldo4;
									elsif respaldo5 > r7 then r7 <= respaldo5;
									elsif respaldo6 > r7 then r7 <= respaldo6;
									elsif data > r7 then r7 <= data; end if;
									salida <= r7;
									cambio_direccion <= '1';
				when "1000" => if respaldo0 > r8 then r8 <= respaldo0;
									elsif respaldo1 > r8 then r8 <= respaldo1;
									elsif respaldo2 > r8 then r8 <= respaldo2; 
									elsif respaldo3 > r8 then r8 <= respaldo3; 
									elsif respaldo4 > r8 then r8 <= respaldo4; 
									elsif respaldo5 > r8 then r8 <= respaldo5;
									elsif respaldo6 > r8 then r8 <= respaldo6; 
									elsif respaldo7 > r8 then r8 <= respaldo7; 
									elsif data > r8 then r8 <= data; end if;
									salida <= r8;
									cambio_direccion <= '1';
				when "1001" => if respaldo0 > r9 then r9 <= respaldo0; 
									elsif respaldo1 > r9 then r9 <= respaldo1; 
									elsif respaldo2 > r9 then r9 <= respaldo2; 
									elsif respaldo3 > r9 then r9 <= respaldo3; 
									elsif respaldo4 > r9 then r9 <= respaldo4; 
									elsif respaldo5 > r9 then r9 <= respaldo5; 
									elsif respaldo6 > r9 then r9 <= respaldo6; 
									elsif respaldo7 > r9 then r9 <= respaldo7; 
									elsif respaldo8 > r9 then r9 <= respaldo8; 
									elsif data > r9 then r9 <= data; end if;
									salida <= r9;
									cambio_direccion <= '1';
				when "1010" => if respaldo0 > r10 then r10 <= respaldo0; 
									elsif respaldo1 > r10 then r10 <= respaldo1; 
									elsif respaldo2 > r10 then r10 <= respaldo2; 
									elsif respaldo3 > r10 then r10 <= respaldo3; 
									elsif respaldo4 > r10 then r10 <= respaldo4; 
									elsif respaldo5 > r10 then r10 <= respaldo5; 
									elsif respaldo6 > r10 then r10 <= respaldo6; 
									elsif respaldo7 > r10 then r10 <= respaldo7; 
									elsif respaldo8 > r10 then r10 <= respaldo8; 
									elsif respaldo9 > r10 then r10 <= respaldo9; 
									elsif data > r10 then r10 <= data; end if;
									salida <= r10;
									cambio_direccion <= '1';
				when "1011" => if respaldo0 > r11 then r11 <= respaldo0; 
									elsif respaldo1 > r11 then r11 <= respaldo1; 
									elsif respaldo2 > r11 then r11 <= respaldo2; 
									elsif respaldo3 > r11 then r11 <= respaldo3; 
									elsif respaldo4 > r11 then r11 <= respaldo4;
									elsif respaldo5 > r11 then r11 <= respaldo5; 
									elsif respaldo6 > r11 then r11 <= respaldo6;
									elsif respaldo7 > r11 then r11 <= respaldo7; 
									elsif respaldo8 > r11 then r11 <= respaldo8; 
									elsif respaldo9 > r11 then r11 <= respaldo9; 
									elsif respaldo10 > r11 then r11 <= respaldo10; 
									elsif data > r11 then r11 <= data; end if;
									salida <= r11;
									cambio_direccion <= '1';
				when "1100" => if respaldo0 > r12 then r12 <= respaldo0; 
									elsif respaldo1 > r12 then r12 <= respaldo1; 
									elsif respaldo2 > r12 then r12 <= respaldo2; 
									elsif respaldo3 > r12 then r12 <= respaldo3; 
									elsif respaldo4 > r12 then r12 <= respaldo4; 
									elsif respaldo5 > r12 then r12 <= respaldo5; 
									elsif respaldo6 > r12 then r12 <= respaldo6; 
									elsif respaldo7 > r12 then r12 <= respaldo7; 
									elsif respaldo8 > r12 then r12 <= respaldo8; 
									elsif respaldo9 > r12 then r12 <= respaldo9; 
									elsif respaldo10 > r12 then r12 <= respaldo10; 
									elsif respaldo11 > r12 then r12 <= respaldo11; 
									elsif data > r12 then r12 <= data; end if;
									salida <= r12;
									cambio_direccion <= '1';
				when "1101" => if respaldo0 > r13 then r13 <= respaldo0; 
									elsif respaldo1 > r13 then r13 <= respaldo1; 
									elsif respaldo2 > r13 then r13 <= respaldo2; 
									elsif respaldo3 > r13 then r13 <= respaldo3; 
									elsif respaldo4 > r13 then r13 <= respaldo4; 
									elsif respaldo5 > r13 then r13 <= respaldo5; 
									elsif respaldo6 > r13 then r13 <= respaldo6; 
									elsif respaldo7 > r13 then r13 <= respaldo7; 
									elsif respaldo8 > r13 then r13 <= respaldo8; 
									elsif respaldo9 > r13 then r13 <= respaldo9; 
									elsif respaldo10 > r13 then r13 <= respaldo10; 
									elsif respaldo11 > r13 then r13 <= respaldo11; 
									elsif respaldo12 > r13 then r13 <= respaldo12;
									elsif data > r13 then r13 <= data; end if;
									salida <= r13;
									cambio_direccion <= '1';
				when "1110" => if respaldo0 > r14 then r14 <= respaldo0; 
									elsif respaldo1 > r14 then r14 <= respaldo1; 
									elsif respaldo2 > r14 then r14 <= respaldo2; 
									elsif respaldo3 > r14 then r14 <= respaldo3; 
									elsif respaldo4 > r14 then r14 <= respaldo4; 
									elsif respaldo5 > r14 then r14 <= respaldo5; 
									elsif respaldo6 > r14 then r14 <= respaldo6; 
									elsif respaldo7 > r14 then r14 <= respaldo7; 
									elsif respaldo8 > r14 then r14 <= respaldo8; 
									elsif respaldo9 > r14 then r14 <= respaldo9; 
									elsif respaldo10 > r14 then r14 <= respaldo10; 
									elsif respaldo11 > r14 then r14 <= respaldo11; 
									elsif respaldo12 > r14 then r14 <= respaldo12; 
									elsif respaldo13 > r14 then r14 <= respaldo13; 
									elsif data > r14 then r14 <= data; end if;
									salida <= r14;
									cambio_direccion <= '1';
				when "1111" => if respaldo0 > r15 then r15 <= respaldo0; 
									elsif respaldo1 > r15 then r15 <= respaldo1; 
									elsif respaldo2 > r15 then r15 <= respaldo2; 
									elsif respaldo3 > r15 then r15 <= respaldo3; 
									elsif respaldo4 > r15 then r15 <= respaldo4; 
									elsif respaldo5 > r15 then r15 <= respaldo5; 
									elsif respaldo6 > r15 then r15 <= respaldo6; 
									elsif respaldo7 > r15 then r15 <= respaldo7; 
									elsif respaldo8 > r15 then r15 <= respaldo8; 
									elsif respaldo9 > r15 then r15 <= respaldo9; 
									elsif respaldo10 > r15 then r15 <= respaldo10; 
									elsif respaldo11 > r15 then r15 <= respaldo11;
									elsif respaldo12 > r15 then r15 <= respaldo12; 
									elsif respaldo13 > r15 then r15 <= respaldo13; 
									elsif respaldo14 > r15 then r15 <= respaldo14; 
									elsif data > r15 then r15 <= data; end if;
									salida <= r15;
									cambio_direccion <= '1';
									cambiar_estado <= '0';
			end case;
		else
			case add is
				when "0000" => q<=r0;
				when "0001" => q<=r1;
				when "0010" => q<=r2;
				when "0011" => q<=r3;
				when "0100" => q<=r4;
				when "0101" => q<=r5;
				when "0110" => q<=r6;
				when "0111" => q<=r7;
				when "1000" => q<=r8;
				when "1001" => q<=r9;
				when "1010" => q<=r10;
				when "1011" => q<=r11;
				when "1100" => q<=r12;
				when "1101" => q<=r13;
				when "1110" => q<=r14;
				when "1111" => q<=r15;
			end case;
		end if;
	end process;
end sol;
